`timescale 1ns / 1ps
/////////////////////////////////////////////////////////////////
// Module Name: four_2_input_or_gate
// Description: Four 2-input OR gate with DELAY configuration parameter
// Parameters: DELAY
/////////////////////////////////////////////////////////////////

module four_2_input_or_gate #(parameter DELAY = 10)(
    input wire a1,b1,a2,b2,a3,b3,a4,b4,
    output wire Y1,Y2,Y3,Y4
    );
    
    or #DELAY (Y1,a1,b1);
    or #DELAY (Y2,a2,b2);
    or #DELAY (Y3,a3,b3);
    or #DELAY (Y4,a4,b4);
    
endmodule
